package apb_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "apb_types.sv"
    `include "apb_item.sv"
    `include "apb_config.sv"

    `include "apb_reg_block.sv"
    `include "apb_reg_adapter.sv"
    `include "apb_sequence.sv"
    `include "apb_slave_sequencer.sv"
    `include "apb_master_sequencer.sv"
    `include "apb_driver.sv"
    `include "apb_master_driver.sv"
    `include "apb_slave_driver.sv"
    `include "apb_monitor.sv"
    `include "apb_slave_agent.sv"
    `include "apb_master_agent.sv"
    `include "apb_predictor.sv"
    `include "apb_scoreboard.sv"

    `include "apb_env.sv"
    `include "apb_test.sv"
endpackage : apb_pkg
